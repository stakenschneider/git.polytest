** Profile: "MAIN-sim"  [ d:\student\myproject\project-main-sim.sim ] 

** Creating circuit file "project-main-sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 16 9.2 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project-MAIN.net" 


.END
